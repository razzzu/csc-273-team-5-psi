module serial_com #(parameter DSIZE=32) (output s_out, r_en
                                input [DSIZE-1:1] rdata,
                                input rempty, rclk, rrst_n);

endmodule
