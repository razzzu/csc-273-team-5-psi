//compile using: vcs -F vcs-psi-compile.txt psi.v

module psi #(parameter DSIZE=32, ASIZE=32) (output s_data, grant, ready,
                                            input [DSIZE-1:0] data,      
                                            input req, pkt_end, p_clk, s_clk, n_rst);

    


endmodule